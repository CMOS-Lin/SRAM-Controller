library verilog;
use verilog.vl_types.all;
entity SRAM_tb is
end SRAM_tb;
